`timescale 1ns / 1ps

module primus_risc_v_top(
  // Input for top module
  input logic clk_i,
  input rst_ni
);

 // logic [31:0]      ir_o          // Instruction register
 // logic [31:0]      npc_o         // Next program counter

 // primus_instruction_fetch a_if (clk_i, rst_ni, pc_i, ir_o, npc_o);
endmodule
